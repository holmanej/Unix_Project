library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library work;
use work.srisc.all;
use work.unix_project.ALL;

entity Unix_Computer is
	port(
		clk			: in  STD_LOGIC
	);
end Unix_Computer;
	
architecture Behavioral of Unix_Computer is

	-- CPU \ IO --
	signal		io_wrData		:	STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal		io_rdData		:	STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal		io_rwAddr		:	STD_LOGIC_VECTOR (3 downto 0) := (others => '0');
	signal		io_wren			:	STD_LOGIC := '0';
	
	-- TEMP GPM --
	signal		guest_pc		:	STD_LOGIC_VECTOR (9 downto 0) := (others => '0');
	signal		guest_insn		:	STD_LOGIC_VECTOR (11 downto 0) := (others => '0');

begin

	CPU: SRISC_CPU port map (
		clk			=> clk,
		reset		=> '0',
		guest_insn	=> guest_insn,
		guest_pc	=> guest_pc,
		io_din		=> io_rdData,
		io_dout		=> io_wrData,
		io_addr		=> io_rwAddr,
		io_wrEn		=> io_wren
	);
	
	IO: IO_Module generic map(x"FF00") port map(
		clk			=> clk,
		cpu_din		=> io_wrData,
		cpu_addr	=> io_rwAddr,
		cpu_wren	=> io_wren,
		cpu_dout	=> io_rdData
	);
	
	GPM: InsnRAM_12bit generic map(10) port map(
		clk			=> clk,
		reset		=> '0',
		-- --
		wrAddr		=> "00000000000",
		wrData		=> x"00",
		wren		=> '0',
		-- --
		rdAddr		=> guest_pc,
		rdData		=> guest_insn
	);

end Behavioral;